module and_32bit(
  input [31:0] a,
  input [31:0] b,
  output [31:0] result
);

  and a0(result[0], a[0], b[0]);
  and a1(result[1], a[1], b[1]);
  and a2(result[2], a[2], b[2]);
  and a3(result[3], a[3], b[3]);
  and a4(result[4], a[4], b[4]);
  and a5(result[5], a[5], b[5]);
  and a6(result[6], a[6], b[6]);
  and a7(result[7], a[7], b[7]);
  and a8(result[8], a[8], b[8]);
  and a9(result[9], a[9], b[9]);
  and a10(result[10], a[10], b[10]);
  and a11(result[11], a[11], b[11]);
  and a12(result[12], a[12], b[12]);
  and a13(result[13], a[13], b[13]);
  and a14(result[14], a[14], b[14]);
  and a15(result[15], a[15], b[15]);
  and a16(result[16], a[16], b[16]);
  and a17(result[17], a[17], b[17]);
  and a18(result[18], a[18], b[18]);
  and a19(result[19], a[19], b[19]);
  and a20(result[20], a[20], b[20]);
  and a21(result[21], a[21], b[21]);
  and a22(result[22], a[22], b[22]);
  and a23(result[23], a[23], b[23]);
  and a24(result[24], a[24], b[24]);
  and a25(result[25], a[25], b[25]);
  and a26(result[26], a[26], b[26]);
  and a27(result[27], a[27], b[27]);
  and a28(result[28], a[28], b[28]);
  and a29(result[29], a[29], b[29]);
  and a30(result[30], a[30], b[30]);
  and a31(result[31], a[31], b[31]);

endmodule
